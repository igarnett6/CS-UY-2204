

module clock_calculator (KEYINPOUT, DIGITENTERED,ENTER,
           ADD, SUB, MUL, DIV, CLEAR, EXP, 
           ADDITION, SUBTRACTION, MULTIPLICATION, DIVISION, EXPONENT,
           AN7, AN6, AN5, AN4, AN3, AN2, AN1, AN0,
           SEGA, SEGB, SEGC, SEGD, SEGE, SEGF, SEGG,
           SETSECOND, SETMINUTE, SETHOUR, SETB, SHOWTIME, 
           TIMERSTARTS, PAUSETIMER, CONTINUETIMER, RESETa, CLK100MHZ,
           ONEHERTZOUT, MODETIMER, MODECLOCK,
           SBUS6, SBUS5, SBUS4, SBUS3, SBUS2, SBUS1, SBUS0, DCDEN7, DCDEN6, DCDEN5, DCDEN4, DCDEN3, DCDEN2, DCDEN1, DCDEN0,
           STREGVAL) ;
         
      
         
///////////////////////////////////////////////////////////////// 
//              Module Declarations Start Below
/////////////////////////////////////////////////////////////////         
         
input DIGITENTERED, ENTER, ADD, SUB, MUL, DIV, CLEAR, EXP, CLK100MHZ ;
inout [7:0] KEYINPOUT ;
output AN7, AN6, AN5, AN4, AN3, AN2, AN1, AN0,SEGA, SEGB, SEGC, SEGD, SEGE, SEGF, SEGG ; 
output ADDITION, SUBTRACTION, MULTIPLICATION, DIVISION, EXPONENT ;
output [4:0] STREGVAL ;

wire signed [15:0] D ;
wire R15, R14, R13, R12, R11, R10, R9, R8, R7, R6, R5, R4, R3, R2, R1, R0 ;
wire [3:0] KEYVAL ;
wire OPRENTERED ;
reg signed [15:0] C ;
reg ADDOP, SUBOP, MULOP, DIVOP, EXPOP ;
reg [3:0] STREG ;
reg signed [7:0] A, B ;
reg ERROR ;
integer i ;
wire RST = 0 ;
wire CLK1HZ, CLK800HZ, CLK100HZ, CLK4HZ ;
reg AE7, AE6, AE5, AE4, AE3, AE2, AE1, AE0 ;
wire OVF ;

//////////////////////////////////////////////////////////////////
//clock declarations start below
/////////////////////////////////////////////////////////////////
input SETSECOND, SETMINUTE, SETHOUR, SHOWTIME, TIMERSTARTS, PAUSETIMER, CONTINUETIMER, RESETa;
input [7:0] SETB;
output ONEHERTZOUT, MODETIMER, MODECLOCK;
output DCDEN7, DCDEN6, DCDEN5, DCDEN4, DCDEN3, DCDEN2, DCDEN1, DCDEN0, SBUS6, SBUS5, SBUS4, SBUS3, SBUS2, SBUS1, SBUS0;

reg [7:0] T;
integer setTime;
integer hoursl, hoursr, secondsl, secondsr, minutesl, minutesr, centisecondsl, centisecondsr;
integer thoursl, thoursr, tsecondsl, tsecondsr, tminutesl, tminutesr, tcentisecondsl, tcentisecondsr;
reg [7:0] H, S ,M, CS;
reg clk, tim;
reg timerON, clockON;

///////////////////////////////////////////////////////////////// 
//             Module Description Starts Below
/////////////////////////////////////////////////////////////////


// Constants are names below

   parameter [4:0] RESET = 5'b00000,
                   S1 = 5'b00001,
                   S2 = 5'b00010,
                   S3 = 5'b00011,
                   S4 = 5'b00100,
                   S5 = 5'b00101,
                   S6 = 5'b00110,
                   S7 = 5'b00111,
                   S8 = 5'b01000,
                   S9 = 5'b01001,
                   S10 = 5'b01010,
                   S11 = 5'b01011,
                   S12 = 5'b01100,
                   S13 = 5'b01101,
                   S14 = 5'b01110,
                   S15 = 5'b01111,
                   S16 = 5'b10000,
                   S17 = 5'b10001,
                   S18 = 5'b10010,
                   S19 = 5'b10011,
                   S20 = 5'b10100,
                   S21 = 5'b10101;
                
                
                                
// Data Unit and Control descriptions start below

// Instantiate the Frequency Divider in the Data Unit
   FREQDIV freq_divider (.ONEHUNDREDMEGAHERTZ(CLK100MHZ), .RESET(RST), 
                         .ONEHERTZ(CLK1HZ), .EIGHTHUNDREDHERTZ(CLK800HZ), .ONEHUNDREDHERTZ(CLK100HZ), .FOURHERTZ(CLK4HZ)) ;
 
 // Instantiate the Key Pad Pmod Controller in the Data Unit
    PmodKEYPAD KeyPad_ctrl (.clk(CLK100MHZ), .JA(KEYINPOUT), .Keypadout(KEYVAL)) ;
   

// Instantiate the ALU Block in the Data Unit
   alu alu_1 (.R15(D[15]), .R14(D[14]), .R13(D[13]), .R12(D[12]), .R11(D[11]), .R10(D[10]), .R9(D[9]), .R8(D[8]),
                         .R7(D[7]), .R6(D[6]), .R5(D[5]), .R4(D[4]), .R3(D[3]), .R2(D[2]), .R1(D[1]), .R0(D[0]), .OVF(OVF), 
                         .K7(A[7]), .K6(A[6]), .K5(A[5]), .K4(A[4]), .K3(A[3]), .K2(A[2]), .K1(A[1]), .K0(A[0]),
                         .M7(B[7]), .M6(B[6]), .M5(B[5]), .M4(B[4]), .M3(B[3]), .M2(B[2]), .M1(B[1]), .M0(B[0]),
                         .ADD(ADDOP), .SUB(SUBOP), .MUL(MULOP), .DIV(DIVOP), .EXP(EXPOP)); 
                         

// Instantiate the 7-Segment Controller in the Data Unit
   ssdCtrl seven_segment_ctrl(.AN7(AN7), .AN6(AN6), .AN5(AN5), .AN4(AN4), .AN3(AN3), .AN2(AN2), .AN1(AN1), .AN0(AN0),
                              .SEGA(SEGA), .SEGB(SEGB), .SEGC(SEGC), .SEGD(SEGD), .SEGE(SEGE), .SEGF(SEGF), .SEGG(SEGG),
                              .CLK100MHZ(CLK100MHZ), .RST(RST), .Err (ERROR),
                              .DIN31(R15), .DIN30(R14), .DIN29(R13), .DIN28(R12), .DIN27(R11), .DIN26(R10), .DIN25(R9), .DIN24(R8), 
                              .DIN23(R7), .DIN22(R6), .DIN21(R5), .DIN20(R4), .DIN19(R3), .DIN18(R2), .DIN17(R1), .DIN16(R0), 
                              .DIN15(B[7]), .DIN14(B[6]), .DIN13(B[5]), .DIN12(B[4]), .DIN11(B[3]), .DIN10(B[2]), .DIN9(B[1]), .DIN8(B[0]), 
                              .DIN7(A[7]), .DIN6(A[6]), .DIN5(A[5]), .DIN4(A[4]), .DIN3(A[3]), .DIN2(A[2]), .DIN1(A[1]), .DIN0(A[0]),
                              .AE7(AE7), .AE6(AE6), .AE5(AE5), .AE4(AE4), .AE3(AE3), .AE2(AE2), .AE1(AE1), .AE0(AE0)) ;
          

// Data Unit circuits
        
    assign OPRENTERED = (ADD | SUB | MUL | DIV | EXP) ;   
  
           
 // Data and Control Unit circuits described together below  
               
   always @ (posedge CLK100HZ) begin
    
        if (clockON == 1) begin // Clock test
            if (centisecondsr == 9) begin
                centisecondsr = 0;
                if (centisecondsl == 9) begin
                    centisecondsl = 0;
                    if (secondsr == 9) begin
                        secondsr = 0;
                        if (secondsl == 5) begin
                            secondsl = 0;
                            if (minutesr == 9) begin
                                minutesr = 0;
                                if (minutesl == 5) begin
                                    minutesl = 0;
                                    if (hoursr == 9) begin
                                        hoursr = 0;
                                            hoursl = hoursl + 1;
                                    end
                                    else if (hoursr == 3 && hoursl == 2) begin
                                        hoursr = 0;
                                        hoursl = 0;
                                    end
                                    else begin
                                        hoursr = hoursr + 1;
                                    end
                                end
                                else begin
                                    minutesl = minutesl + 1;
                                end
                            end
                            else begin
                                minutesr = minutesr + 1;
                            end
                        end
                        else begin
                            secondsl = secondsl + 1;
                        end
                    end
                    else begin
                        secondsr = secondsr + 1;
                    end
                end
                else begin
                    centisecondsl = centisecondsl + 1;
                end
            end
            else begin
                centisecondsr = centisecondsr + 1;
            end
        end
    
        if (timerON == 1) begin // timer test
                if (tcentisecondsr == 9) begin
                    tcentisecondsr = 0;
                    if (tcentisecondsl == 9) begin
                        tcentisecondsl = 0;
                        if (tsecondsr == 9) begin
                            tsecondsr = 0;
                            if (tsecondsl == 5) begin
                                tsecondsl = 0;
                                if (tminutesr == 9) begin
                                    tminutesr = 0;
                                    if (tminutesl == 5) begin
                                        tminutesl = 0;
                                        if (thoursr == 9) begin
                                            thoursr = 0;
                                                thoursl = thoursl + 1;
                                        end
                                        else if (thoursr == 3 && thoursl == 2) begin
                                            thoursr = 0;
                                            thoursl = 0;
                                        end
                                        else begin
                                            thoursr = hoursr + 1;
                                        end
                                    end
                                    else begin
                                        tminutesl = tminutesl + 1;
                                    end
                                end
                                else begin
                                    tminutesr = tminutesr + 1;
                                end
                            end
                            else begin
                                tsecondsl = tsecondsl + 1;
                            end
                        end
                        else begin
                            tsecondsr = tsecondsr + 1;
                        end
                    end
                    else begin
                        tcentisecondsl = tcentisecondsl + 1;
                    end
                end
                else begin
                    tcentisecondsr = tcentisecondsr + 1;
                end
            end
        
    
        
        
       case (STREG)
          RESET : begin H <= 8'd0 ; M <= 8'd0 ; S <= 8'd0 ; CS <= 8'd0 ; 
                        tim <= 0;
                        clk = 0;
                        clockON <= 0;
                        timerON <= 0;
                        hoursl = 0;
                        minutesl = 0;
                        secondsl = 0;
                        centisecondsl = 0;
                        thoursl = 0;
                        tminutesl = 0;
                        tsecondsl = 0;
                        tcentisecondsl = 0;
                        hoursr = 0;
                        minutesr = 0;
                        secondsr = 0;
                        centisecondsr = 0;
                        thoursr = 0;
                        tminutesr = 0;
                        tsecondsr = 0;
                        tcentisecondsr = 0;
                        
                        AE7<= 0 ; AE6<= 0 ; AE5<= 0 ; AE4<=0 ; AE3<= 0 ; AE2<= 0 ; AE1<= 0 ; AE0<= 0 ; 
                        
                         if (RESETa) STREG <= RESET ;
                         else if (SETSECOND) STREG <= S1 ; 
                         else if (SETMINUTE) STREG <= S2 ;
                         else if (SETHOUR) STREG <= S3 ;
                         else if (SHOWTIME) STREG <= S4 ;
                  end
  
          S1 : begin i <= SETB ; AE2 <= 0 ; AE3 <= 0; 
                     secondsl = i/10;
                     secondsr = i%10;
                     S[3:0] <= secondsr;
                     S[7:4] <= secondsl;
                     if (RESETa) STREG <= RESET ;
                     else if (SETSECOND) STREG <= S1 ; 
                     else if (SETMINUTE) STREG <= S2 ;
                     else if (SETHOUR) STREG <= S3 ; // not in state diagram but this is more helpful for user
                     else if (SHOWTIME) STREG <= S4 ;
               end
                
          S2 : begin i <= SETB ; AE4 <= 0 ; AE5 <= 0;
                    minutesl <= i/10;
                    minutesr <= i%10;
                    M[7:4] <= minutesl;
                    M[3:0] <= minutesr;
                    if (RESETa) STREG <= RESET ;
                    else if (SETSECOND) STREG <= S1 ; // not in state diagram but this is more helpful for user
                    else if (SETMINUTE) STREG <= S2 ;
                    else if (SETHOUR) STREG <= S3 ;
                    else if (SHOWTIME) STREG <= S4 ;
               end           
          
          S3 : begin i <= SETB ; AE6 <= 0 ; AE7 <= 0;
                    hoursl = i/10;
                    hoursr = i%10;
                    H[7:4] <= hoursl;
                    H[3:0] <= hoursr;
                    if (RESETa) STREG <= RESET ;
                    else if (SETSECOND) STREG <= S1 ; // not in state diagram but this is more helpful for user
                    else if (SETMINUTE) STREG <= S2 ; // not in state diagram but this is more helpful for user
                    else if (SETHOUR) STREG <= S3 ;
                    else if (SHOWTIME) STREG <= S4 ;
               end
          
          S4 : begin clockON <= 1;
               AE7<= 0 ; AE6<= 0 ; AE5<= 0 ; AE4<=0 ; AE3<= 0 ; AE2<= 0 ; AE1<= 0 ; AE0<= 0 ; 
               clk <= 1;
               H[7:4] <= hoursl;
               H[3:0] <= hoursr;
               M[7:4] <= minutesl;
               M[3:0] <= minutesr;
               S[7:4] <= secondsl;
               S[3:0] <= secondsr;
               CS[7:4] <= centisecondsl;
               CS[3:0] <= centisecondsr;
               if (RESETa) STREG <= RESET ;
               else if (SETSECOND) STREG <= S1 ;
               else if (SETMINUTE) STREG <= S2 ;
               else if (SETHOUR) STREG <= S3 ;
               else if (TIMERSTARTS) STREG <= S5 ;
               else if (PAUSETIMER) STREG <= S6 ;
               else if (CONTINUETIMER) STREG <= S7 ; 
               end
                
                
          S5 : begin CS[7:0] <= SETB ; 
                   AE7<= 0 ; AE6<= 0 ; AE5<= 0 ; AE4<=0 ; AE3<= 0 ; AE2<= 0 ; AE1<= 0 ; AE0<= 0 ; 
                   timerON <= 1;
                   tim <=1;
                   clk <= 0;
                   H[7:4] <= thoursl;
                   H[3:0] <= thoursr;
                   M[7:4] <= tminutesl;
                   M[3:0] <= tminutesr;
                   S[7:4] <= tsecondsl;
                   S[3:0] <= tsecondsr;
                   CS[7:4] <= tcentisecondsl;
                   CS[3:0] <= tcentisecondsr;
                   if (RESETa) STREG <= RESET ;
                   else if (SHOWTIME) STREG <= S4 ;
                   else if (TIMERSTARTS) STREG <= S5 ;
                   else if (PAUSETIMER) STREG <= S6 ;                   
               end
          
          S6 : begin CS[7:0] <= SETB ;
                   AE7<= 0 ; AE6<= 0 ; AE5<= 0 ; AE4<=0 ; AE3<= 0 ; AE2<= 0 ; AE1<= 0 ; AE0<= 0 ; 
                   timerON <= 0;
                   tim <=0;
                   clk <= 0;
                   if (RESETa) STREG <= RESET ;
                   else if (SHOWTIME) STREG <= S4 ;
                   else if (PAUSETIMER) STREG <= S6 ;   
                   else if (CONTINUETIMER) STREG <= S7 ;                  
               end
               
          S7 : begin CS[7:0] <= SETB ; 
                   AE7<= 0 ; AE6<= 0 ; AE5<= 0 ; AE4<=0 ; AE3<= 0 ; AE2<= 0 ; AE1<= 0 ; AE0<= 0 ; 
                   timerON <= 1;
                   tim <= 1;
                   clk <= 0;
                   H[7:4] <= thoursl;
                   H[3:0] <= thoursr;
                   M[7:4] <= tminutesl;
                   M[3:0] <= tminutesr;
                   S[7:4] <= tsecondsl;
                   S[3:0] <= tsecondsr;
                   CS[7:4] <= tcentisecondsl;
                   CS[3:0] <= tcentisecondsr;
                   if (RESETa) STREG <= RESET ;
                   else if (SHOWTIME) STREG <= S4 ;
                   else if (CONTINUETIMER) STREG <= S7 ; 
               end
    
    
    
    //START OF CALCULATOR STATES
    
    
    
 
          S8 : begin C <= 16'd0 ; A <= 8'd0 ; B <= 8'd0 ; 
                        ADDOP <= 0 ; SUBOP <= 0 ; MULOP <= 0 ; DIVOP <= 0 ; EXPOP <= 0 ; ERROR <= 0 ;
                        AE7<= 1 ; AE6<= 1 ; AE5<= 1 ; AE4<=1 ; AE3<= 1 ; AE2<= 1 ; AE1<= 1 ; AE0<= 1 ; 
                         if (CLEAR) STREG <= RESET ;
                             else if (DIGITENTERED) STREG <= S9 ; 
                  end
  
          S9 : begin A[3:0] <= KEYVAL ; AE0 <= 0 ; 
                     if (CLEAR) STREG <= RESET ;
                          else if (~DIGITENTERED) STREG <= S10 ;
               end
                
          S10 :  if (CLEAR) STREG <= RESET ;
                    else if (DIGITENTERED) STREG <= S11 ;
                             else if (OPRENTERED)          
                                      begin
                                         STREG <= S13 ; 
                                         if (ADD) begin  ADDOP <= 1 ; SUBOP <= 0 ; MULOP <= 0 ; DIVOP <= 0 ; EXPOP <= 0 ; end
                                             else if (SUB) begin ADDOP <= 0 ; SUBOP <= 1 ; MULOP <= 0 ; DIVOP <= 0 ; EXPOP <= 0 ; end
                                                     else if (MUL) begin ADDOP <= 0 ; SUBOP <= 0 ; MULOP <= 1 ; DIVOP <= 0 ; EXPOP <= 0 ; end
                                                             else if (DIV) begin ADDOP <= 0 ; SUBOP <= 0 ; MULOP <= 0 ; DIVOP <= 1 ; EXPOP <= 0 ; end
                                                                      else if (EXP) begin ADDOP <= 0 ; SUBOP <= 0 ; MULOP <= 0 ; DIVOP <= 0 ; EXPOP <= 1 ; end 
                                     end 
          
          S11 : begin if (A[3:0] != 0) begin A[7:4] <= A[3:0] ; AE1 <= 0 ; end
                     if (CLEAR) STREG <= RESET ;
                         else if (~DIGITENTERED) STREG <= S12 ; 
               end      
          
          S12 : begin A[3:0] <= KEYVAL ; 
                     if (CLEAR) STREG <= RESET ;
                         else if (OPRENTERED)
                                  begin
                                       STREG <= S13 ; 
                                       if (ADD) begin  ADDOP <= 1 ; SUBOP <= 0 ; MULOP <= 0 ; DIVOP <= 0 ; EXPOP <= 0 ; end
                                           else if (SUB) begin ADDOP <= 0 ; SUBOP <= 1 ; MULOP <= 0 ; DIVOP <= 0 ; EXPOP <= 0 ; end
                                                else if (MUL) begin ADDOP <= 0 ; SUBOP <= 0 ; MULOP <= 1 ; DIVOP <= 0 ; EXPOP <= 0 ; end
                                                   else if (DIV) begin ADDOP <= 0 ; SUBOP <= 0 ; MULOP <= 0 ; DIVOP <= 1 ; EXPOP <= 0 ; end
                                                            else if (EXP) begin ADDOP <= 0 ; SUBOP <= 0 ; MULOP <= 0 ; DIVOP <= 0 ; EXPOP <= 1 ; end 
                                 end 
                end
                
          S13 : begin
                    if (ADD) begin  ADDOP <= 1 ; SUBOP <= 0 ; MULOP <= 0 ; DIVOP <= 0 ; EXPOP <= 0 ; end
                       else if (SUB) begin ADDOP <= 0 ; SUBOP <= 1 ; MULOP <= 0 ; DIVOP <= 0 ; EXPOP <= 0 ; end
                                else if (MUL) begin ADDOP <= 0 ; SUBOP <= 0 ; MULOP <= 1 ; DIVOP <= 0 ; EXPOP <= 0 ; end
                                        else if (DIV) begin ADDOP <= 0 ; SUBOP <= 0 ; MULOP <= 0 ; DIVOP <= 1 ; EXPOP <= 0 ; end 
                                                 else if (EXP) begin ADDOP <= 0 ; SUBOP <= 0 ; MULOP <= 0 ; DIVOP <= 0 ; EXPOP <= 1 ; end
                  if (CLEAR) STREG <= RESET ;
                  else if (DIGITENTERED) STREG <= S14 ; 
               end
          
          S14 : begin B[3:0] <= KEYVAL ; AE2 <= 0 ; 
                     if (CLEAR) STREG <= RESET ;
                         else if (~DIGITENTERED) STREG <= S15 ;
               end
               
          S15 : if (CLEAR) STREG <= RESET ;
                  else if (DIGITENTERED) STREG <= S16 ;
                           else if (ENTER)STREG <= S10 ;       
          
          S16 : begin if (B[3:0] != 0) begin B[7:4] <= B[3:0] ; AE3 <= 0 ; end 
                     if (CLEAR) STREG <= RESET ;
                         if (~DIGITENTERED) STREG <= S17 ;
                end
          
          S17 :  begin B[3:0] <= KEYVAL ; 
                      if (CLEAR) STREG <= RESET ;
                          else if (ENTER) STREG <= S18 ;
               end
          
          S18 : begin if (((B == 8'd0) & DIVOP) | ((B[7] == 1) & EXPOP) | (OVF)) ERROR <= 1 ;
                      else C <= D ;
                      if (CLEAR) STREG <= RESET ;
                         else STREG <= S19 ; 
                end
                
          S19 :  begin if ((C[3:0] != 0) | (C[7:4] != 0) | (C[11:8] != 0)| (C[15:12] != 0))  AE4<= 0;
                       if ((C[7:4] != 0) | (C[11:8] != 0)| (C[15:12] != 0)) AE5 <=0;
                       if ((C[11:8] != 0) | (C[15:12] != 0)) AE6 <=0;
                       if (C[15:12] != 0) AE7<= 0;
                       if (CLEAR) STREG <= RESET ;
                         else if (DIGITENTERED) STREG <= S20 ; 
                 end           
          
          S20 : begin C <= 16'd0 ; A <= 8'd0 ; B <= 8'd0 ; 
                     ADDOP <= 0 ; SUBOP <= 0 ; MULOP <= 0 ; DIVOP <= 0 ; EXPOP <= 0 ;ERROR <= 0 ;
                     AE7<= 1 ; AE6<= 1 ; AE5<= 1 ; AE4<=1 ; AE3<= 1 ; AE2<= 1 ; AE1<= 1 ; AE0<= 1 ;
                     if (CLEAR == 1) STREG <= RESET ;
                        else STREG <= S21 ;
                end                               
          
          S21 : begin if (KEYVAL != 0) begin A[3:0] <= KEYVAL ; AE0 <= 0 ; end
                      if (CLEAR) STREG <= RESET ;
                          else if (~DIGITENTERED) STREG <= S10 ;
                end
          
          default STREG <= RESET ;
        endcase
     end                       
       
       
// Data Unit circuits below
                                                  
//  The ADDITION, SUBTRACTION, MULTIPLICATION and DIVISION LED light ouputs receive their values from their registers

       assign {R15, R14, R13, R12, R11, R10, R9, R8, R7, R6, R5, R4, R3, R2, R1, R0} = C ;
       assign ADDITION = ADDOP;
       assign SUBTRACTION = SUBOP ;
       assign MULTIPLICATION = MULOP ;
       assign DIVISION = DIVOP ;
       assign EXPONENT = EXPOP ;
       assign STREGVAL = STREG ;
   
   
/////////////////////////////////////////////////////////////////


endmodule